module ALU( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222613.2]
  input  [3:0]  io_fn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222616.4]
  input  [31:0] io_in2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222616.4]
  input  [31:0] io_in1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222616.4]
  output [31:0] io_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222616.4]
  output [31:0] io_adder_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222616.4]
  output        io_cmp_out // @[:freechips.rocketchip.system.DefaultRV32Config.fir@222616.4]
);
  wire [31:0] _T_1; // @[ALU.scala 62:35:freechips.rocketchip.system.DefaultRV32Config.fir@222622.4]
  wire [31:0] in2_inv; // @[ALU.scala 62:20:freechips.rocketchip.system.DefaultRV32Config.fir@222623.4]
  wire [31:0] in1_xor_in2; // @[ALU.scala 63:28:freechips.rocketchip.system.DefaultRV32Config.fir@222624.4]
  wire [31:0] _T_3; // @[ALU.scala 64:26:freechips.rocketchip.system.DefaultRV32Config.fir@222626.4]
  wire [31:0] _GEN_0; // @[ALU.scala 64:36:freechips.rocketchip.system.DefaultRV32Config.fir@222628.4]
  wire  _T_9; // @[ALU.scala 68:24:freechips.rocketchip.system.DefaultRV32Config.fir@222633.4]
  wire  _T_14; // @[ALU.scala 69:8:freechips.rocketchip.system.DefaultRV32Config.fir@222638.4]
  wire  slt; // @[ALU.scala 68:8:freechips.rocketchip.system.DefaultRV32Config.fir@222639.4]
  wire  _T_17; // @[ALU.scala 44:26:freechips.rocketchip.system.DefaultRV32Config.fir@222642.4]
  wire  _T_18; // @[ALU.scala 70:68:freechips.rocketchip.system.DefaultRV32Config.fir@222643.4]
  wire  _T_19; // @[ALU.scala 70:41:freechips.rocketchip.system.DefaultRV32Config.fir@222644.4]
  wire [4:0] shamt; // @[ALU.scala 74:28:freechips.rocketchip.system.DefaultRV32Config.fir@222647.4]
  wire  _T_21; // @[ALU.scala 82:24:freechips.rocketchip.system.DefaultRV32Config.fir@222648.4]
  wire  _T_22; // @[ALU.scala 82:44:freechips.rocketchip.system.DefaultRV32Config.fir@222649.4]
  wire  _T_23; // @[ALU.scala 82:35:freechips.rocketchip.system.DefaultRV32Config.fir@222650.4]
  wire [31:0] _T_27; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222654.4]
  wire [31:0] _T_29; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222656.4]
  wire [31:0] _T_31; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222658.4]
  wire [31:0] _T_32; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222659.4]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222664.4]
  wire [31:0] _T_37; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222664.4]
  wire [31:0] _T_39; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222666.4]
  wire [31:0] _T_41; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222668.4]
  wire [31:0] _T_42; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222669.4]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222674.4]
  wire [31:0] _T_47; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222674.4]
  wire [31:0] _T_49; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222676.4]
  wire [31:0] _T_51; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222678.4]
  wire [31:0] _T_52; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222679.4]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222684.4]
  wire [31:0] _T_57; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222684.4]
  wire [31:0] _T_59; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222686.4]
  wire [31:0] _T_61; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222688.4]
  wire [31:0] _T_62; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222689.4]
  wire [31:0] _GEN_4; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222694.4]
  wire [31:0] _T_67; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222694.4]
  wire [31:0] _T_69; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222696.4]
  wire [31:0] _T_71; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222698.4]
  wire [31:0] _T_72; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222699.4]
  wire [31:0] shin; // @[ALU.scala 82:17:freechips.rocketchip.system.DefaultRV32Config.fir@222700.4]
  wire  _T_75; // @[ALU.scala 83:35:freechips.rocketchip.system.DefaultRV32Config.fir@222703.4]
  wire [32:0] _T_77; // @[ALU.scala 83:57:freechips.rocketchip.system.DefaultRV32Config.fir@222705.4]
  wire [32:0] _T_78; // @[ALU.scala 83:64:freechips.rocketchip.system.DefaultRV32Config.fir@222706.4]
  wire [31:0] shout_r; // @[ALU.scala 83:73:freechips.rocketchip.system.DefaultRV32Config.fir@222707.4]
  wire [31:0] _T_82; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222711.4]
  wire [31:0] _T_84; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222713.4]
  wire [31:0] _T_86; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222715.4]
  wire [31:0] _T_87; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222716.4]
  wire [31:0] _GEN_5; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222721.4]
  wire [31:0] _T_92; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222721.4]
  wire [31:0] _T_94; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222723.4]
  wire [31:0] _T_96; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222725.4]
  wire [31:0] _T_97; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222726.4]
  wire [31:0] _GEN_6; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222731.4]
  wire [31:0] _T_102; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222731.4]
  wire [31:0] _T_104; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222733.4]
  wire [31:0] _T_106; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222735.4]
  wire [31:0] _T_107; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222736.4]
  wire [31:0] _GEN_7; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222741.4]
  wire [31:0] _T_112; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222741.4]
  wire [31:0] _T_114; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222743.4]
  wire [31:0] _T_116; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222745.4]
  wire [31:0] _T_117; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222746.4]
  wire [31:0] _GEN_8; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222751.4]
  wire [31:0] _T_122; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222751.4]
  wire [31:0] _T_124; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222753.4]
  wire [31:0] _T_126; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222755.4]
  wire [31:0] shout_l; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222756.4]
  wire [31:0] _T_130; // @[ALU.scala 85:18:freechips.rocketchip.system.DefaultRV32Config.fir@222760.4]
  wire  _T_131; // @[ALU.scala 86:25:freechips.rocketchip.system.DefaultRV32Config.fir@222761.4]
  wire [31:0] _T_132; // @[ALU.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@222762.4]
  wire [31:0] shout; // @[ALU.scala 85:74:freechips.rocketchip.system.DefaultRV32Config.fir@222763.4]
  wire  _T_133; // @[ALU.scala 89:25:freechips.rocketchip.system.DefaultRV32Config.fir@222764.4]
  wire  _T_134; // @[ALU.scala 89:45:freechips.rocketchip.system.DefaultRV32Config.fir@222765.4]
  wire  _T_135; // @[ALU.scala 89:36:freechips.rocketchip.system.DefaultRV32Config.fir@222766.4]
  wire [31:0] _T_136; // @[ALU.scala 89:18:freechips.rocketchip.system.DefaultRV32Config.fir@222767.4]
  wire  _T_138; // @[ALU.scala 90:44:freechips.rocketchip.system.DefaultRV32Config.fir@222769.4]
  wire  _T_139; // @[ALU.scala 90:35:freechips.rocketchip.system.DefaultRV32Config.fir@222770.4]
  wire [31:0] _T_140; // @[ALU.scala 90:63:freechips.rocketchip.system.DefaultRV32Config.fir@222771.4]
  wire [31:0] _T_141; // @[ALU.scala 90:18:freechips.rocketchip.system.DefaultRV32Config.fir@222772.4]
  wire [31:0] logic_; // @[ALU.scala 89:78:freechips.rocketchip.system.DefaultRV32Config.fir@222773.4]
  wire  _T_142; // @[ALU.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@222774.4]
  wire  _T_143; // @[ALU.scala 91:35:freechips.rocketchip.system.DefaultRV32Config.fir@222775.4]
  wire [31:0] _GEN_9; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@222776.4]
  wire [31:0] _T_144; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@222776.4]
  wire [31:0] shift_logic; // @[ALU.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@222777.4]
  wire  _T_145; // @[ALU.scala 92:23:freechips.rocketchip.system.DefaultRV32Config.fir@222778.4]
  wire  _T_146; // @[ALU.scala 92:43:freechips.rocketchip.system.DefaultRV32Config.fir@222779.4]
  wire  _T_147; // @[ALU.scala 92:34:freechips.rocketchip.system.DefaultRV32Config.fir@222780.4]
  assign _T_1 = ~io_in2; // @[ALU.scala 62:35:freechips.rocketchip.system.DefaultRV32Config.fir@222622.4]
  assign in2_inv = io_fn[3] ? _T_1 : io_in2; // @[ALU.scala 62:20:freechips.rocketchip.system.DefaultRV32Config.fir@222623.4]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 63:28:freechips.rocketchip.system.DefaultRV32Config.fir@222624.4]
  assign _T_3 = io_in1 + in2_inv; // @[ALU.scala 64:26:freechips.rocketchip.system.DefaultRV32Config.fir@222626.4]
  assign _GEN_0 = {{31'd0}, io_fn[3]}; // @[ALU.scala 64:36:freechips.rocketchip.system.DefaultRV32Config.fir@222628.4]
  assign _T_9 = io_in1[31] == io_in2[31]; // @[ALU.scala 68:24:freechips.rocketchip.system.DefaultRV32Config.fir@222633.4]
  assign _T_14 = io_fn[1] ? io_in2[31] : io_in1[31]; // @[ALU.scala 69:8:freechips.rocketchip.system.DefaultRV32Config.fir@222638.4]
  assign slt = _T_9 ? io_adder_out[31] : _T_14; // @[ALU.scala 68:8:freechips.rocketchip.system.DefaultRV32Config.fir@222639.4]
  assign _T_17 = ~io_fn[3]; // @[ALU.scala 44:26:freechips.rocketchip.system.DefaultRV32Config.fir@222642.4]
  assign _T_18 = in1_xor_in2 == 32'h0; // @[ALU.scala 70:68:freechips.rocketchip.system.DefaultRV32Config.fir@222643.4]
  assign _T_19 = _T_17 ? _T_18 : slt; // @[ALU.scala 70:41:freechips.rocketchip.system.DefaultRV32Config.fir@222644.4]
  assign shamt = io_in2[4:0]; // @[ALU.scala 74:28:freechips.rocketchip.system.DefaultRV32Config.fir@222647.4]
  assign _T_21 = io_fn == 4'h5; // @[ALU.scala 82:24:freechips.rocketchip.system.DefaultRV32Config.fir@222648.4]
  assign _T_22 = io_fn == 4'hb; // @[ALU.scala 82:44:freechips.rocketchip.system.DefaultRV32Config.fir@222649.4]
  assign _T_23 = _T_21 | _T_22; // @[ALU.scala 82:35:freechips.rocketchip.system.DefaultRV32Config.fir@222650.4]
  assign _T_27 = {{16'd0}, io_in1[31:16]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222654.4]
  assign _T_29 = {io_in1[15:0], 16'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222656.4]
  assign _T_31 = _T_29 & 32'hffff0000; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222658.4]
  assign _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222659.4]
  assign _GEN_1 = {{8'd0}, _T_32[31:8]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222664.4]
  assign _T_37 = _GEN_1 & 32'hff00ff; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222664.4]
  assign _T_39 = {_T_32[23:0], 8'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222666.4]
  assign _T_41 = _T_39 & 32'hff00ff00; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222668.4]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222669.4]
  assign _GEN_2 = {{4'd0}, _T_42[31:4]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222674.4]
  assign _T_47 = _GEN_2 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222674.4]
  assign _T_49 = {_T_42[27:0], 4'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222676.4]
  assign _T_51 = _T_49 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222678.4]
  assign _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222679.4]
  assign _GEN_3 = {{2'd0}, _T_52[31:2]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222684.4]
  assign _T_57 = _GEN_3 & 32'h33333333; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222684.4]
  assign _T_59 = {_T_52[29:0], 2'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222686.4]
  assign _T_61 = _T_59 & 32'hcccccccc; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222688.4]
  assign _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222689.4]
  assign _GEN_4 = {{1'd0}, _T_62[31:1]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222694.4]
  assign _T_67 = _GEN_4 & 32'h55555555; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222694.4]
  assign _T_69 = {_T_62[30:0], 1'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222696.4]
  assign _T_71 = _T_69 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222698.4]
  assign _T_72 = _T_67 | _T_71; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222699.4]
  assign shin = _T_23 ? io_in1 : _T_72; // @[ALU.scala 82:17:freechips.rocketchip.system.DefaultRV32Config.fir@222700.4]
  assign _T_75 = io_fn[3] & shin[31]; // @[ALU.scala 83:35:freechips.rocketchip.system.DefaultRV32Config.fir@222703.4]
  assign _T_77 = {_T_75,shin}; // @[ALU.scala 83:57:freechips.rocketchip.system.DefaultRV32Config.fir@222705.4]
  assign _T_78 = $signed(_T_77) >>> shamt; // @[ALU.scala 83:64:freechips.rocketchip.system.DefaultRV32Config.fir@222706.4]
  assign shout_r = _T_78[31:0]; // @[ALU.scala 83:73:freechips.rocketchip.system.DefaultRV32Config.fir@222707.4]
  assign _T_82 = {{16'd0}, shout_r[31:16]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222711.4]
  assign _T_84 = {shout_r[15:0], 16'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222713.4]
  assign _T_86 = _T_84 & 32'hffff0000; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222715.4]
  assign _T_87 = _T_82 | _T_86; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222716.4]
  assign _GEN_5 = {{8'd0}, _T_87[31:8]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222721.4]
  assign _T_92 = _GEN_5 & 32'hff00ff; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222721.4]
  assign _T_94 = {_T_87[23:0], 8'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222723.4]
  assign _T_96 = _T_94 & 32'hff00ff00; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222725.4]
  assign _T_97 = _T_92 | _T_96; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222726.4]
  assign _GEN_6 = {{4'd0}, _T_97[31:4]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222731.4]
  assign _T_102 = _GEN_6 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222731.4]
  assign _T_104 = {_T_97[27:0], 4'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222733.4]
  assign _T_106 = _T_104 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222735.4]
  assign _T_107 = _T_102 | _T_106; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222736.4]
  assign _GEN_7 = {{2'd0}, _T_107[31:2]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222741.4]
  assign _T_112 = _GEN_7 & 32'h33333333; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222741.4]
  assign _T_114 = {_T_107[29:0], 2'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222743.4]
  assign _T_116 = _T_114 & 32'hcccccccc; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222745.4]
  assign _T_117 = _T_112 | _T_116; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222746.4]
  assign _GEN_8 = {{1'd0}, _T_117[31:1]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222751.4]
  assign _T_122 = _GEN_8 & 32'h55555555; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@222751.4]
  assign _T_124 = {_T_117[30:0], 1'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@222753.4]
  assign _T_126 = _T_124 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@222755.4]
  assign shout_l = _T_122 | _T_126; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@222756.4]
  assign _T_130 = _T_23 ? shout_r : 32'h0; // @[ALU.scala 85:18:freechips.rocketchip.system.DefaultRV32Config.fir@222760.4]
  assign _T_131 = io_fn == 4'h1; // @[ALU.scala 86:25:freechips.rocketchip.system.DefaultRV32Config.fir@222761.4]
  assign _T_132 = _T_131 ? shout_l : 32'h0; // @[ALU.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@222762.4]
  assign shout = _T_130 | _T_132; // @[ALU.scala 85:74:freechips.rocketchip.system.DefaultRV32Config.fir@222763.4]
  assign _T_133 = io_fn == 4'h4; // @[ALU.scala 89:25:freechips.rocketchip.system.DefaultRV32Config.fir@222764.4]
  assign _T_134 = io_fn == 4'h6; // @[ALU.scala 89:45:freechips.rocketchip.system.DefaultRV32Config.fir@222765.4]
  assign _T_135 = _T_133 | _T_134; // @[ALU.scala 89:36:freechips.rocketchip.system.DefaultRV32Config.fir@222766.4]
  assign _T_136 = _T_135 ? in1_xor_in2 : 32'h0; // @[ALU.scala 89:18:freechips.rocketchip.system.DefaultRV32Config.fir@222767.4]
  assign _T_138 = io_fn == 4'h7; // @[ALU.scala 90:44:freechips.rocketchip.system.DefaultRV32Config.fir@222769.4]
  assign _T_139 = _T_134 | _T_138; // @[ALU.scala 90:35:freechips.rocketchip.system.DefaultRV32Config.fir@222770.4]
  assign _T_140 = io_in1 & io_in2; // @[ALU.scala 90:63:freechips.rocketchip.system.DefaultRV32Config.fir@222771.4]
  assign _T_141 = _T_139 ? _T_140 : 32'h0; // @[ALU.scala 90:18:freechips.rocketchip.system.DefaultRV32Config.fir@222772.4]
  assign logic_ = _T_136 | _T_141; // @[ALU.scala 89:78:freechips.rocketchip.system.DefaultRV32Config.fir@222773.4]
  assign _T_142 = io_fn >= 4'hc; // @[ALU.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@222774.4]
  assign _T_143 = _T_142 & slt; // @[ALU.scala 91:35:freechips.rocketchip.system.DefaultRV32Config.fir@222775.4]
  assign _GEN_9 = {{31'd0}, _T_143}; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@222776.4]
  assign _T_144 = _GEN_9 | logic_; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@222776.4]
  assign shift_logic = _T_144 | shout; // @[ALU.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@222777.4]
  assign _T_145 = io_fn == 4'h1; // @[ALU.scala 92:23:freechips.rocketchip.system.DefaultRV32Config.fir@222778.4]
  assign _T_146 = io_fn == 4'ha; // @[ALU.scala 92:43:freechips.rocketchip.system.DefaultRV32Config.fir@222779.4]
  assign _T_147 = _T_145 | _T_146; // @[ALU.scala 92:34:freechips.rocketchip.system.DefaultRV32Config.fir@222780.4]
  assign io_out = _T_147 ? io_adder_out : shift_logic; // @[ALU.scala 94:10:freechips.rocketchip.system.DefaultRV32Config.fir@222782.4]
  assign io_adder_out = _T_3 + _GEN_0; // @[ALU.scala 64:16:freechips.rocketchip.system.DefaultRV32Config.fir@222630.4]
  assign io_cmp_out = io_fn[0] ^ _T_19; // @[ALU.scala 70:14:freechips.rocketchip.system.DefaultRV32Config.fir@222646.4]
endmodule
